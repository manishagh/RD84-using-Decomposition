library IEEE;
use IEEE.std_logic_1164.all;


entity G1 is 
 	port(
 x: in STD_LOGIC_VECTOR(0 to 2);
 y: out STD_LOGIC_VECTOR(0 to 1) );
 end G1;
 
architecture G1 of G1 is 
 begin
 	 with x select 
 		    y <= 
"00" when "000",
	
"01" when "100",
	
"01" when "010",
	
"10" when "110",
	
"01" when "001",
	
"10" when "101",
	
"10" when "011",
	
"11" when "111",
	
"--" when others; 
 end G1;
 
 library IEEE;
use IEEE.std_logic_1164.all;


entity G2 is 
 	port(
 x: in STD_LOGIC_VECTOR(0 to 2);
 y: out STD_LOGIC_VECTOR(0 to 1) );
 end G2;
 
architecture G2 of G2 is 
 begin
 	 with x select 
 		    y <= 
"00" when "000",
	
"01" when "001",
	
"01" when "100",
	
"10" when "101",
	
"01" when "010",
	
"10" when "011",
	
"10" when "110",
	
"11" when "111",
	
"--" when others; 
 end G2;
 
library IEEE;
use IEEE.std_logic_1164.all;


entity G3 is 
 	port(
 x: in STD_LOGIC_VECTOR(0 to 2);
 y: out STD_LOGIC_VECTOR(0 to 1) );
 end G3;
 
architecture G3 of G3 is 
 begin
 	 with x select 
 		    y <= 
"00" when "000",
	
"01" when "001",
	
"01" when "100",
	
"10" when "101",
	
"01" when "010",
	
"10" when "011",
	
"10" when "110",
	
"11" when "111",
	
"--" when others; 
 end G3;
 
 library IEEE;
use IEEE.std_logic_1164.all;


entity H_rd84 is 
 	port(
 x: in STD_LOGIC_VECTOR(0 to 4);
 y: out STD_LOGIC_VECTOR(0 to 3) );
 end H_rd84;
 
architecture H_rd84 of H_rd84 is 
 begin
 	 with x select 
 		    y <= 
"0000" when "00000",
	
"0100" when "00001",
	
"0100" when "00100",
	
"1000" when "00101",
	
"1000" when "01000",
	
"1100" when "01001",
	
"1000" when "10000",
	
"1100" when "10100",
	
"0001" when "11000",
	
"1000" when "00010",
	
"1100" when "00110",
	
"0001" when "01010",
	
"1100" when "10001",
	
"0001" when "10101",
	
"0101" when "11001",
	
"1100" when "01100",
	
"0001" when "01101",
	
"0101" when "11100",
	
"0101" when "01110",
	
"1001" when "11101",
	
"0001" when "10010",
	
"0101" when "10110",
	
"1001" when "11010",
	
"1101" when "11110",
	
"1100" when "00011",
	
"0001" when "00111",
	
"0101" when "01011",
	
"1001" when "01111",
	
"0101" when "10011",
	
"1001" when "10111",
	
"1101" when "11011",
	
"0010" when "11111",
	
"----" when others; 
 end H_rd84;
 
library IEEE;
use IEEE.std_logic_1164.all;


entity rd84 is 
 	port(
 x: in STD_LOGIC_VECTOR(0 to 7);
 y: out STD_LOGIC_VECTOR(0 to 3) );
 end rd84;
 
 architecture rd84 of rd84 is
 component G1 
      port(
  x: in STD_LOGIC_VECTOR(0 to 2);
  y: out STD_LOGIC_VECTOR(0 to 1) );
      end component;
      
     component G2 
           port(
       x: in STD_LOGIC_VECTOR(0 to 2);
       y: out STD_LOGIC_VECTOR(0 to 1) );
     end component; 
     
     component G3 
          port(
      x: in STD_LOGIC_VECTOR(0 to 2);
      y: out STD_LOGIC_VECTOR(0 to 1) );
     end component;
     
     component H_rd84 
           port(
      x: in STD_LOGIC_VECTOR(0 to 4);
      y: out STD_LOGIC_VECTOR(0 to 3) );
           end component;
 signal temp1, temp2, temp3 : std_logic_vector(0 to 1);
 signal a,b: std_logic_vector(0 to 2);
 signal c: std_logic_vector(0 to 4);
 begin 
 --d<=x(0)&x(1)&x(2);
 uut1: G1 port map (x(0 to 2),temp1);
 a<=temp1&x(3);
 uut2: G2 port map (a,temp2);
 b<=temp2&x(5);
 uut3: G3 port map (b,temp3);
 c<= x(4)&temp3&x(6)&x(7);
 uut4: H_rd84 port map(c,y);
 end;
 --end rd84;

library ieee;
use ieee.std_logic_1164.all;

entity TbTt is
 end TbTt;

 architecture mytest of tbtt is

signal x: std_logic_vector (0 to 7);
 signal y: std_logic_vector (0 to 3); 
type test_vector is record
	x: std_logic_vector (0 to 7);
 	 y:  std_logic_vector (0 to 3);
 end record;
 
type test_vector_array is array (natural range <>) of test_vector;
	constant test_vectors: test_vector_array := (

	(x => "00000000", y => "0000"),

	(x => "10000000", y => "0100"),

	(x => "00000100", y => "0100"),

	(x => "10000100", y => "1000"),

	(x => "00010000", y => "0100"),

	(x => "10010000", y => "1000"),

	(x => "00010100", y => "1000"),

	(x => "10010100", y => "1100"),

	(x => "01000000", y => "0100"),

	(x => "11000000", y => "1000"),

	(x => "01000100", y => "1000"),

	(x => "11000100", y => "1100"),

	(x => "01010000", y => "1000"),

	(x => "11010000", y => "1100"),

	(x => "01010100", y => "1100"),

	(x => "11010100", y => "0001"),

	(x => "00000010", y => "0100"),

	(x => "10000010", y => "1000"),

	(x => "00000110", y => "1000"),

	(x => "10000110", y => "1100"),

	(x => "00010010", y => "1000"),

	(x => "10010010", y => "1100"),

	(x => "00010110", y => "1100"),

	(x => "10010110", y => "0001"),

	(x => "01000010", y => "1000"),

	(x => "11000010", y => "1100"),

	(x => "01000110", y => "1100"),

	(x => "11000110", y => "0001"),

	(x => "01010010", y => "1100"),

	(x => "11010010", y => "0001"),

	(x => "01010110", y => "0001"),

	(x => "11010110", y => "0101"),

	(x => "00001000", y => "0100"),

	(x => "10001000", y => "1000"),

	(x => "00001100", y => "1000"),

	(x => "10001100", y => "1100"),

	(x => "00011000", y => "1000"),

	(x => "10011000", y => "1100"),

	(x => "00011100", y => "1100"),

	(x => "10011100", y => "0001"),

	(x => "01001000", y => "1000"),

	(x => "11001000", y => "1100"),

	(x => "01001100", y => "1100"),

	(x => "11001100", y => "0001"),

	(x => "01011000", y => "1100"),

	(x => "11011000", y => "0001"),

	(x => "01011100", y => "0001"),

	(x => "11011100", y => "0101"),

	(x => "00001010", y => "1000"),

	(x => "10001010", y => "1100"),

	(x => "00001110", y => "1100"),

	(x => "10001110", y => "0001"),

	(x => "00011010", y => "1100"),

	(x => "10011010", y => "0001"),

	(x => "00011110", y => "0001"),

	(x => "10011110", y => "0101"),

	(x => "01001010", y => "1100"),

	(x => "11001010", y => "0001"),

	(x => "01001110", y => "0001"),

	(x => "11001110", y => "0101"),

	(x => "01011010", y => "0001"),

	(x => "11011010", y => "0101"),

	(x => "01011110", y => "0101"),

	(x => "11011110", y => "1001"),

	(x => "00100000", y => "0100"),

	(x => "10100000", y => "1000"),

	(x => "00100100", y => "1000"),

	(x => "10100100", y => "1100"),

	(x => "00110000", y => "1000"),

	(x => "10110000", y => "1100"),

	(x => "00110100", y => "1100"),

	(x => "10110100", y => "0001"),

	(x => "01100000", y => "1000"),

	(x => "11100000", y => "1100"),

	(x => "01100100", y => "1100"),

	(x => "11100100", y => "0001"),

	(x => "01110000", y => "1100"),

	(x => "11110000", y => "0001"),

	(x => "01110100", y => "0001"),

	(x => "11110100", y => "0101"),

	(x => "00100010", y => "1000"),

	(x => "10100010", y => "1100"),

	(x => "00100110", y => "1100"),

	(x => "10100110", y => "0001"),

	(x => "00110010", y => "1100"),

	(x => "10110010", y => "0001"),

	(x => "00110110", y => "0001"),

	(x => "10110110", y => "0101"),

	(x => "01100010", y => "1100"),

	(x => "11100010", y => "0001"),

	(x => "01100110", y => "0001"),

	(x => "11100110", y => "0101"),

	(x => "01110010", y => "0001"),

	(x => "11110010", y => "0101"),

	(x => "01110110", y => "0101"),

	(x => "11110110", y => "1001"),

	(x => "00101000", y => "1000"),

	(x => "10101000", y => "1100"),

	(x => "00101100", y => "1100"),

	(x => "10101100", y => "0001"),

	(x => "00111000", y => "1100"),

	(x => "10111000", y => "0001"),

	(x => "00111100", y => "0001"),

	(x => "10111100", y => "0101"),

	(x => "01101000", y => "1100"),

	(x => "11101000", y => "0001"),

	(x => "01101100", y => "0001"),

	(x => "11101100", y => "0101"),

	(x => "01111000", y => "0001"),

	(x => "11111000", y => "0101"),

	(x => "01111100", y => "0101"),

	(x => "11111100", y => "1001"),

	(x => "00101010", y => "1100"),

	(x => "10101010", y => "0001"),

	(x => "00101110", y => "0001"),

	(x => "10101110", y => "0101"),

	(x => "00111010", y => "0001"),

	(x => "10111010", y => "0101"),

	(x => "00111110", y => "0101"),

	(x => "10111110", y => "1001"),

	(x => "01101010", y => "0001"),

	(x => "11101010", y => "0101"),

	(x => "01101110", y => "0101"),

	(x => "11101110", y => "1001"),

	(x => "01111010", y => "0101"),

	(x => "11111010", y => "1001"),

	(x => "01111110", y => "1001"),

	(x => "11111110", y => "1101"),

	(x => "00000001", y => "0100"),

	(x => "10000001", y => "1000"),

	(x => "00000101", y => "1000"),

	(x => "10000101", y => "1100"),

	(x => "00010001", y => "1000"),

	(x => "10010001", y => "1100"),

	(x => "00010101", y => "1100"),

	(x => "10010101", y => "0001"),

	(x => "01000001", y => "1000"),

	(x => "11000001", y => "1100"),

	(x => "01000101", y => "1100"),

	(x => "11000101", y => "0001"),

	(x => "01010001", y => "1100"),

	(x => "11010001", y => "0001"),

	(x => "01010101", y => "0001"),

	(x => "11010101", y => "0101"),

	(x => "00000011", y => "1000"),

	(x => "10000011", y => "1100"),

	(x => "00000111", y => "1100"),

	(x => "10000111", y => "0001"),

	(x => "00010011", y => "1100"),

	(x => "10010011", y => "0001"),

	(x => "00010111", y => "0001"),

	(x => "10010111", y => "0101"),

	(x => "01000011", y => "1100"),

	(x => "11000011", y => "0001"),

	(x => "01000111", y => "0001"),

	(x => "11000111", y => "0101"),

	(x => "01010011", y => "0001"),

	(x => "11010011", y => "0101"),

	(x => "01010111", y => "0101"),

	(x => "11010111", y => "1001"),

	(x => "00001001", y => "1000"),

	(x => "10001001", y => "1100"),

	(x => "00001101", y => "1100"),

	(x => "10001101", y => "0001"),

	(x => "00011001", y => "1100"),

	(x => "10011001", y => "0001"),

	(x => "00011101", y => "0001"),

	(x => "10011101", y => "0101"),

	(x => "01001001", y => "1100"),

	(x => "11001001", y => "0001"),

	(x => "01001101", y => "0001"),

	(x => "11001101", y => "0101"),

	(x => "01011001", y => "0001"),

	(x => "11011001", y => "0101"),

	(x => "01011101", y => "0101"),

	(x => "11011101", y => "1001"),

	(x => "00001011", y => "1100"),

	(x => "10001011", y => "0001"),

	(x => "00001111", y => "0001"),

	(x => "10001111", y => "0101"),

	(x => "00011011", y => "0001"),

	(x => "10011011", y => "0101"),

	(x => "00011111", y => "0101"),

	(x => "10011111", y => "1001"),

	(x => "01001011", y => "0001"),

	(x => "11001011", y => "0101"),

	(x => "01001111", y => "0101"),

	(x => "11001111", y => "1001"),

	(x => "01011011", y => "0101"),

	(x => "11011011", y => "1001"),

	(x => "01011111", y => "1001"),

	(x => "11011111", y => "1101"),

	(x => "00100001", y => "1000"),

	(x => "10100001", y => "1100"),

	(x => "00100101", y => "1100"),

	(x => "10100101", y => "0001"),

	(x => "00110001", y => "1100"),

	(x => "10110001", y => "0001"),

	(x => "00110101", y => "0001"),

	(x => "10110101", y => "0101"),

	(x => "01100001", y => "1100"),

	(x => "11100001", y => "0001"),

	(x => "01100101", y => "0001"),

	(x => "11100101", y => "0101"),

	(x => "01110001", y => "0001"),

	(x => "11110001", y => "0101"),

	(x => "01110101", y => "0101"),

	(x => "11110101", y => "1001"),

	(x => "00100011", y => "1100"),

	(x => "10100011", y => "0001"),

	(x => "00100111", y => "0001"),

	(x => "10100111", y => "0101"),

	(x => "00110011", y => "0001"),

	(x => "10110011", y => "0101"),

	(x => "00110111", y => "0101"),

	(x => "10110111", y => "1001"),

	(x => "01100011", y => "0001"),

	(x => "11100011", y => "0101"),

	(x => "01100111", y => "0101"),

	(x => "11100111", y => "1001"),

	(x => "01110011", y => "0101"),

	(x => "11110011", y => "1001"),

	(x => "01110111", y => "1001"),

	(x => "11110111", y => "1101"),

	(x => "00101001", y => "1100"),

	(x => "10101001", y => "0001"),

	(x => "00101101", y => "0001"),

	(x => "10101101", y => "0101"),

	(x => "00111001", y => "0001"),

	(x => "10111001", y => "0101"),

	(x => "00111101", y => "0101"),

	(x => "10111101", y => "1001"),

	(x => "01101001", y => "0001"),

	(x => "11101001", y => "0101"),

	(x => "01101101", y => "0101"),

	(x => "11101101", y => "1001"),

	(x => "01111001", y => "0101"),

	(x => "11111001", y => "1001"),

	(x => "01111101", y => "1001"),

	(x => "11111101", y => "1101"),

	(x => "00101011", y => "0001"),

	(x => "10101011", y => "0101"),

	(x => "00101111", y => "0101"),

	(x => "10101111", y => "1001"),

	(x => "00111011", y => "0101"),

	(x => "10111011", y => "1001"),

	(x => "00111111", y => "1001"),

	(x => "10111111", y => "1101"),

	(x => "01101011", y => "0101"),

	(x => "11101011", y => "1001"),

	(x => "01101111", y => "1001"),

	(x => "11101111", y => "1101"),

	(x => "01111011", y => "1001"),

	(x => "11111011", y => "1101"),

	(x => "01111111", y => "1101"),

	(x => "11111111", y => "0010"));

component rd84 is
	 port(
 x: in STD_LOGIC_VECTOR(0 to 7);
 y: out STD_LOGIC_VECTOR(0 to 3)
);
end component;
 
begin
uut: rd84 port map(x, y);
 	 verify: process  	variable vector: test_vector;  	variable error: boolean:= false;
 	begin 
 	      for i in test_vectors' range loop
	          vector := test_vectors(i); 
      x <= vector.x;  
    wait for 20 ns;

 	        if y /= vector.y then
 		         assert false report"y is wrong value";
error:= true;
end if;
end loop;
assert not error report "Test vectors failed." severity note;
 assert error report "Test vectors passed." severity note;
 wait;
 end process;
end; 
